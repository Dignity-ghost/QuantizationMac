module mac();













endmodule